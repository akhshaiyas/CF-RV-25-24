/*
see LICENSE.iitm
--------------------------------------------------------------------------------------------------
*/
`define number_of_multiplier_stages 4
`define multiplier_latency 5
`define XLEN 64

